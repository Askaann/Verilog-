// verilog code Full Adder
module Full_Adder(A,B,Cin,Sum,Cout);
  input A,B,Cin;
  output Sum,Cout;

  Half_adder
